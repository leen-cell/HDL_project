// adder for four bit number made of four full adders , sums two numbers each made of 4 bits
module Adder (sum,carryout,A,B,c);
//inputs and outputs
input c ;
input[3:0] A,B ;
output carryout;
output [3:0]sum;
wire c1,c2,c3;
 //instantiate four full adders
FA num1 (sum[0],c1,A[0],B[0],c);
FA num2 (sum[1],c2,A[1],B[1],c1);
FA num3 (sum[2],c3,A[2],B[2],c2);
FA num4 (sum[3],carryout,A[3],B[3],c3);
endmodule 